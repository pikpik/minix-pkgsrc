@comment $NetBSD$
${CT_WEBDIR}/system/modules/backend/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/backend/languages/sv/countries.php
${CT_WEBDIR}/system/modules/backend/languages/sv/default.php
${CT_WEBDIR}/system/modules/backend/languages/sv/explain.php
${CT_WEBDIR}/system/modules/backend/languages/sv/languages.php
${CT_WEBDIR}/system/modules/backend/languages/sv/modules.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_article.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_content.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_files.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_form.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_form_field.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_install.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_layout.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_log.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_maintenance.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_member.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_member_group.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_page.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_settings.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_style.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_style_sheet.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_task.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_theme.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_undo.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_user.php
${CT_WEBDIR}/system/modules/backend/languages/sv/tl_user_group.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/calendar/languages/sv/default.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/modules.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/tl_calendar.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/tl_calendar_events.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/tl_user.php
${CT_WEBDIR}/system/modules/calendar/languages/sv/tl_user_group.php
${CT_WEBDIR}/system/modules/comments/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/comments/languages/sv/modules.php
${CT_WEBDIR}/system/modules/comments/languages/sv/tl_comments.php
${CT_WEBDIR}/system/modules/comments/languages/sv/tl_content.php
${CT_WEBDIR}/system/modules/comments/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/faq/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/faq/languages/sv/default.php
${CT_WEBDIR}/system/modules/faq/languages/sv/modules.php
${CT_WEBDIR}/system/modules/faq/languages/sv/tl_faq.php
${CT_WEBDIR}/system/modules/faq/languages/sv/tl_faq_category.php
${CT_WEBDIR}/system/modules/faq/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/frontend/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/frontend/languages/sv/default.php
${CT_WEBDIR}/system/modules/frontend/languages/sv/modules.php
${CT_WEBDIR}/system/modules/listing/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/listing/languages/sv/modules.php
${CT_WEBDIR}/system/modules/listing/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/news/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/news/languages/sv/default.php
${CT_WEBDIR}/system/modules/news/languages/sv/modules.php
${CT_WEBDIR}/system/modules/news/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/news/languages/sv/tl_news.php
${CT_WEBDIR}/system/modules/news/languages/sv/tl_news_archive.php
${CT_WEBDIR}/system/modules/news/languages/sv/tl_news_comments.php
${CT_WEBDIR}/system/modules/news/languages/sv/tl_user.php
${CT_WEBDIR}/system/modules/news/languages/sv/tl_user_group.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/newsletter/languages/sv/default.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/modules.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_member.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_newsletter.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_newsletter_channel.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_newsletter_recipients.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_user.php
${CT_WEBDIR}/system/modules/newsletter/languages/sv/tl_user_group.php
${CT_WEBDIR}/system/modules/registration/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/registration/languages/sv/default.php
${CT_WEBDIR}/system/modules/registration/languages/sv/modules.php
${CT_WEBDIR}/system/modules/registration/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/rep_base/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/rep_base/languages/sv/modules.php
${CT_WEBDIR}/system/modules/rep_base/languages/sv/tl_repository.php
${CT_WEBDIR}/system/modules/rep_base/languages/sv/tl_settings.php
${CT_WEBDIR}/system/modules/rep_client/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/rep_client/languages/sv/modules.php
${CT_WEBDIR}/system/modules/rep_client/languages/sv/tl_repository.php
${CT_WEBDIR}/system/modules/rep_client/languages/sv/tl_settings.php
${CT_WEBDIR}/system/modules/rss_reader/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/rss_reader/languages/sv/modules.php
${CT_WEBDIR}/system/modules/rss_reader/languages/sv/tl_module.php
${CT_WEBDIR}/system/modules/tpl_editor/languages/sv/.htaccess
${CT_WEBDIR}/system/modules/tpl_editor/languages/sv/modules.php
${CT_WEBDIR}/system/modules/tpl_editor/languages/sv/tl_templates.php
