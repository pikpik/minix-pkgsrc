@comment $NetBSD$
${DRUPAL_BASE}/LICENSE.sv.txt
${DRUPAL_BASE}/STATUS.sv.txt
${DRUPAL_BASE}/modules/system/translations/general.sv.po
${DRUPAL_BASE}/modules/system/translations/includes.sv.po
${DRUPAL_BASE}/profiles/default/translations/sv.po
${DRUPAL_BASE}/modules/system/translations/misc.sv.po
${DRUPAL_BASE}/modules/aggregator/translations/modules-aggregator.sv.po
${DRUPAL_BASE}/modules/block/translations/modules-block.sv.po
${DRUPAL_BASE}/modules/blog/translations/modules-blog.sv.po
${DRUPAL_BASE}/modules/blogapi/translations/modules-blogapi.sv.po
${DRUPAL_BASE}/modules/book/translations/modules-book.sv.po
${DRUPAL_BASE}/modules/color/translations/modules-color.sv.po
${DRUPAL_BASE}/modules/comment/translations/modules-comment.sv.po
${DRUPAL_BASE}/modules/contact/translations/modules-contact.sv.po
${DRUPAL_BASE}/modules/dblog/translations/modules-dblog.sv.po
${DRUPAL_BASE}/modules/filter/translations/modules-filter.sv.po
${DRUPAL_BASE}/modules/forum/translations/modules-forum.sv.po
${DRUPAL_BASE}/modules/help/translations/modules-help.sv.po
${DRUPAL_BASE}/modules/locale/translations/modules-locale.sv.po
${DRUPAL_BASE}/modules/menu/translations/modules-menu.sv.po
${DRUPAL_BASE}/modules/node/translations/modules-node.sv.po
${DRUPAL_BASE}/modules/openid/translations/modules-openid.sv.po
${DRUPAL_BASE}/modules/path/translations/modules-path.sv.po
${DRUPAL_BASE}/modules/php/translations/modules-php.sv.po
${DRUPAL_BASE}/modules/ping/translations/modules-ping.sv.po
${DRUPAL_BASE}/modules/poll/translations/modules-poll.sv.po
${DRUPAL_BASE}/modules/profile/translations/modules-profile.sv.po
${DRUPAL_BASE}/modules/search/translations/modules-search.sv.po
${DRUPAL_BASE}/modules/statistics/translations/modules-statistics.sv.po
${DRUPAL_BASE}/modules/syslog/translations/modules-syslog.sv.po
${DRUPAL_BASE}/modules/system/translations/modules-system.sv.po
${DRUPAL_BASE}/modules/taxonomy/translations/modules-taxonomy.sv.po
${DRUPAL_BASE}/modules/throttle/translations/modules-throttle.sv.po
${DRUPAL_BASE}/modules/tracker/translations/modules-tracker.sv.po
${DRUPAL_BASE}/modules/translation/translations/modules-translation.sv.po
${DRUPAL_BASE}/modules/trigger/translations/modules-trigger.sv.po
${DRUPAL_BASE}/modules/update/translations/modules-update.sv.po
${DRUPAL_BASE}/modules/upload/translations/modules-upload.sv.po
${DRUPAL_BASE}/modules/user/translations/modules-user.sv.po
${DRUPAL_BASE}/themes/chameleon/translations/themes-chameleon.sv.po
${DRUPAL_BASE}/themes/garland/translations/themes-garland.sv.po
${DRUPAL_BASE}/themes/pushbutton/translations/themes-pushbutton.sv.po
